LIBRARY ieee;
USE ieee.STD_LOGIC_1164.all; 

ENTITY DESLOCADOR_L IS
	PORT(
		CK, CLR, SET: IN STD_LOGIC;
		DIR, ESQ: IN STD_LOGIC; -- CHAVE DIRE��O DO DESLOCAMENTO S1 DIR E S2 LEFT
		D: OUT STD_LOGIC_VECTOR (0 TO 7) -- DESLOCAMENTO 
);
END DESLOCADOR_L;

  
ARCHITECTURE DESLOCADOR_F OF DESLOCADOR_L IS
	COMPONENT ffd is
  	port (ck, clr, set, d : in  std_logic;
              q : out std_logic);
	END COMPONENT FFD;

	
	COMPONENT MUX_2_ENTSEL IS
	PORT(
		A00, A01, A10, A11: IN STD_LOGIC; --ENTRADAS
		S0, S1: IN STD_LOGIC; --ENTRADA SELE��O
		Q: OUT STD_LOGIC --SAIDA
	);
	END COMPONENT MUX_2_ENTSEL;
	
	SIGNAL Q : STD_LOGIC_VECTOR(0 TO 7);
	SIGNAL SM: STD_LOGIC_VECTOR(0 TO 7); --SAIDA MUX

BEGIN	
	--COMPONENTE REG_MUX_0
	MUX0 : MUX_2_ENTSEL PORT MAP(Q(0), Q(7), Q(1),Q(0), DIR, ESQ, SM(0));
	FFD0 : ffd PORT MAP(CK, CLR, SET, SM(0), Q(0));

	--COMPONENTE REG_MUX_1
	MUX1 : MUX_2_ENTSEL PORT MAP(Q(1), Q(0), Q(2),Q(1), DIR, ESQ, SM(1));
	FFD1 : ffd PORT MAP(CK, CLR, '1', SM(1), Q(1));

	--COMPONENTE REG_MUX_2
	MUX2 : MUX_2_ENTSEL PORT MAP(Q(2), Q(1), Q(3),Q(2), DIR, ESQ, SM(2));
	FFD2 : ffd PORT MAP(CK, CLR, '1', SM(2), Q(2));

	--COMPONENTE REG_MUX_3
	MUX3 : MUX_2_ENTSEL PORT MAP(Q(3), Q(2), Q(4),Q(3), DIR, ESQ, SM(3));
	FFD3 : ffd PORT MAP(CK, CLR, '1', SM(3), Q(3));

	--COMPONENTE REG_MUX_4
	MUX4 : MUX_2_ENTSEL PORT MAP(Q(4), Q(3), Q(5),Q(4), DIR, ESQ, SM(4));
	FFD4 : ffd PORT MAP(CK, CLR, '1', SM(4), Q(4));

	--COMPONENTE REG_MUX_5
	MUX5 : MUX_2_ENTSEL PORT MAP(Q(5), Q(4), Q(6),Q(5), DIR, ESQ, SM(5));
	FFD5 : ffd PORT MAP(CK, CLR, '1', SM(5), Q(5));

	--COMPONENTE REG_MUX_6
	MUX6 : MUX_2_ENTSEL PORT MAP(Q(6), Q(5), Q(7),Q(6), DIR, ESQ, SM(6));
	FFD6 : ffd PORT MAP(CK, CLR, '1', SM(6), Q(6));

	--COMPONENTE REG_MUX_7
	MUX7 : MUX_2_ENTSEL PORT MAP(Q(7), Q(6), Q(0),Q(7), DIR, ESQ, SM(7));
	FFD7 : ffd PORT MAP(CK, CLR, '1', SM(7), Q(7));

	D(0) <= Q(0);
	D(1) <= Q(1);
	D(2) <= Q(2);
	D(3) <= Q(3);
	D(4) <= Q(4);
	D(5) <= Q(5);
	D(6) <= Q(6);
	D(7) <= Q(7);

END DESLOCADOR_F;
