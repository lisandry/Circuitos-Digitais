LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY COMPARADOR_4BIT is
	Port(
		A, B: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		EQ, GT, LT: OUT STD_LOGIC
);
END ENTITY COMPARADOR_4BIT;


ARCHITECTURE COMPARADOR_4BIT OF COMPARADOR_4BIT IS  

	COMPONENT COMPARADOR_1BIT is
	Port(
		A, B: IN STD_LOGIC;
		EQ, GT, LT: OUT STD_LOGIC
	);
	END COMPONENT COMPARADOR_1BIT;
	
	SIGNAL EQ3, GT3, LT3, EQ2, GT2, LT2, EQ1, GT1, LT1, EQ0, GT0, LT0 : STD_LOGIC;

BEGIN
C3 : COMPARADOR_1BIT PORT MAP (A(3), B(3), EQ3, GT3, LT3);
C2 : COMPARADOR_1BIT PORT MAP (A(2), B(2), EQ2, GT2, LT2);
C1 : COMPARADOR_1BIT PORT MAP (A(1), B(1), EQ1, GT1, LT1);
C0 : COMPARADOR_1BIT PORT MAP (A(0), B(0), EQ0, GT0, LT0);

EQ <= EQ3 AND EQ2 AND EQ1 AND EQ0;
GT <= GT3 OR GT2 OR GT1 OR GT0;
LT <= NOT(EQ3 AND EQ2 AND EQ1 AND EQ0) AND NOT(GT3 OR GT2 OR GT1 OR GT0);

END ARCHITECTURE COMPARADOR_4BIT;
