LIBRARY ieee;
USE ieee.STD_LOGIC_1164.all;

ENTITY MUX_2_ENTSEL IS
	PORT(
		A00, A01, A10, A11: IN STD_LOGIC; --ENTRADAS
		S0, S1: IN STD_LOGIC; --ENTRADA SELE��O
		Q: OUT STD_LOGIC --SAIDA
);
END MUX_2_ENTSEL;

ARCHITECTURE MUX_2_ENTSEL OF MUX_2_ENTSEL IS
	SIGNAL A_00, A_01, A_10, A_11: STD_LOGIC;
	
BEGIN

	A_00 <= (NOT(S1) AND NOT(S0)) AND A00;
	A_01 <= (NOT(S1) AND S0) AND A01;
	A_10 <= (S1 AND NOT(S0)) AND A10;
	A_11 <= (S1 AND S0) AND A11;

	Q <= A_00 OR A_01 OR A_10 OR A_11;

END ARCHITECTURE;


