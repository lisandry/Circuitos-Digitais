LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY BLOCO_RC IS
	PORT(
		CLR_R, LOAD_R, LOAD_C, CLK: IN STD_LOGIC;
		Y_IN, C: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		Y_OUT: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		PROD_YC: OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
);
END BLOCO_RC;

ARCHITECTURE BLOCO_RC OF BLOCO_RC IS

	COMPONENT REG_C IS
	PORT(
		LOAD_C, CLK: IN STD_LOGIC;
		D: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		S: OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
	);
	END COMPONENT REG_C;

	COMPONENT REG_Y IS
	PORT(
		CLR_R, LOAD_R, CLK: IN STD_LOGIC;
		D: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		S: OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
	);
	END COMPONENT REG_Y;

	COMPONENT MULTIPLICADOR_4BITS IS
	PORT(
		A, B: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		R: OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
	);
	END COMPONENT MULTIPLICADOR_4BITS;

	SIGNAL C_AUX, Y_AUX: STD_LOGIC_VECTOR(3 DOWNTO 0);

BEGIN

REGC: REG_C PORT MAP (LOAD_C, CLK, C, C_AUX);
REGY: REG_Y PORT MAP (CLR_R ,LOAD_R, CLK, Y_IN, Y_AUX);

Y_OUT <= Y_AUX;

MULT: MULTIPLICADOR_4BITS PORT MAP (C_AUX, Y_AUX, PROD_YC);

END ARCHITECTURE BLOCO_RC;
