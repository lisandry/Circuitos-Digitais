LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY COMPARADOR_1BIT is
	Port(
		A, B: IN STD_LOGIC;
		EQ, GT, LT: OUT STD_LOGIC
);
END ENTITY COMPARADOR_1BIT;
	
ARCHITECTURE COMPARADOR_1BIT OF COMPARADOR_1BIT IS
BEGIN

LT <= NOT(A) AND B;
GT <= A AND NOT(B);
EQ <= (NOT(A) AND NOT(B)) OR (A AND B);

END ARCHITECTURE COMPARADOR_1BIT;