LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY COD_2X4 IS
	PORT(
		EN: IN STD_LOGIC;
		S1, S0: IN STD_LOGIC;
		Q3, Q2, Q1, Q0: OUT STD_LOGIC
);
END COD_2X4;
		
ARCHITECTURE CODIFICADOR_2X4 OF COD_2X4 IS

BEGIN
	Q3 <= EN AND S1 AND S0;
	Q2 <= EN AND S1 AND (NOT(S0));
	Q1 <= EN AND (NOT(S1)) AND S0;
	Q0 <= EN AND (NOT(S1)) AND (NOT(S0));

END ARCHITECTURE;
	
