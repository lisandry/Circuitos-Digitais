LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY MULTIPLICADOR_4BITS IS
	PORT(
		A, B: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		R: OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
);
END MULTIPLICADOR_4BITS;

ARCHITECTURE MULTIPLICADOR OF MULTIPLICADOR_4BITS IS
	COMPONENT Somador_Completo is
        PORT(
        	A_SC, B_SC, CI_SC: IN STD_LOGIC;
        	S_SC, CO_SC: OUT STD_LOGIC
        );
    	END COMPONENT;

	--SIGNAL ENTRADAS SOMADOR 0
	SIGNAL A00, A01, A02, A03: STD_LOGIC;
	SIGNAL B00, B01, B02, B03: STD_LOGIC;
	SIGNAL CA00, CA01, CA02, CA03: STD_LOGIC;

	--SIGNAL ENTRADAS SOMADOR 1
	SIGNAL A10, A11, A12, A13: STD_LOGIC;
	SIGNAL B10, B11, B12, B13, B14, B15: STD_LOGIC;
	SIGNAL CA10, CA11, CA12, CA13, CA14: STD_LOGIC;

	--SIGNAL ENTRADAS SOMADOR 2
	SIGNAL A20, A21, A22, A23: STD_LOGIC;
	SIGNAL B20, B21, B22, B23, B24, B25, B26: STD_LOGIC;
	SIGNAL CA20, CA21, CA22, CA23, CA24, CA25: STD_LOGIC;

	--SIGNAL COUT DOS SOMADORES
	SIGNAL CA_OUT0, CA_OUT1, CA_OUT2: STD_LOGIC;

	--SIGNAL SAIDA SOMADOR 0
	SIGNAL S00, S01, S02, S03, S04: STD_LOGIC;

	--SIGNAL SAIDA SOMADOR 1
	SIGNAL S10, S11, S12, S13, S14, S15: STD_LOGIC;

	--SIGNAL SAIDA SOMADOR 2
	SIGNAL S20, S21, S22, S23, S24, S25, S26: STD_LOGIC;




BEGIN

-- ENTRADAS SOMADOR 0
A00 <= A(0) AND B(0);
A01 <= A(1) AND B(0);
A02 <= A(2) AND B(0);
A03 <= A(3) AND B(0);


B00 <= A(0) AND B(1);
B01 <= A(1) AND B(1);
B02 <= A(2) AND B(1);
B03 <= A(3) AND B(1);

--SOMADOR 0
S_AB00: Somador_Completo PORT MAP(A00,'0', '0',S00 , CA00);
S_AB01: Somador_Completo PORT MAP(A01,B00, CA00,S01 ,CA01);
S_AB02: Somador_Completo PORT MAP(A02,B01, CA01,S02 ,CA02);
S_AB03: Somador_Completo PORT MAP(A03,B02, CA02,S03 ,CA03);
S_AB04: Somador_Completo PORT MAP('0',B03, CA03,S04 ,CA_OUT0);

-- ENTRADAS SOMADOR 1
A10 <= A(0) AND B(2);
A11 <= A(1) AND B(2);
A12 <= A(2) AND B(2);
A13 <= A(3) AND B(2);


B10 <= S00;
B11 <= S01;
B12 <= S02;
B13 <= S03;
B14 <= S04;
B15 <= CA_OUT0;

--SOMADOR 1
S_AB10: Somador_Completo PORT MAP('0',B10, '0',  S10 ,CA10);
S_AB11: Somador_Completo PORT MAP('0',B11, CA10, S11 ,CA11);
S_AB12: Somador_Completo PORT MAP(A10,B12, CA11, S12 ,CA12);
S_AB13: Somador_Completo PORT MAP(A11,B13, CA12, S13 ,CA13);
S_AB14: Somador_Completo PORT MAP(A12,B14, CA13, S14 ,CA14);
S_AB15: Somador_Completo PORT MAP(A13,B15, CA14, S15 ,CA_OUT1);

-- ENTRADAS SOMADOR 2
A20 <= A(0) AND B(3);
A21 <= A(1) AND B(3);
A22 <= A(2) AND B(3);
A23 <= A(3) AND B(3);


B20 <= S10;
B21 <= S11;
B22 <= S12;
B23 <= S13;
B24 <= S14;
B25 <= S15;
B26 <= CA_OUT1;

--SOMADOR 2
S_AB20: Somador_Completo PORT MAP('0',B20, '0',  S20 ,CA20);
S_AB21: Somador_Completo PORT MAP('0',B21, CA20, S21 ,CA21);
S_AB22: Somador_Completo PORT MAP('0',B22, CA21, S22 ,CA22);
S_AB23: Somador_Completo PORT MAP(A20,B23, CA22, S23 ,CA23);
S_AB24: Somador_Completo PORT MAP(A21,B24, CA23 ,S24 ,CA24);
S_AB25: Somador_Completo PORT MAP(A22,B25, CA24, S25 ,CA25);
S_AB26: Somador_Completo PORT MAP(A23,B26, CA25, S26 ,CA_OUT2);


--RESULTADO
R(0) <= S20;
R(1) <= S21;
R(2) <= S22;
R(3) <= S23;
R(4) <= S24;
R(5) <= S25;
R(6) <= S26;
R(7) <= CA_OUT2;

END ARCHITECTURE MULTIPLICADOR;